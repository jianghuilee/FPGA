module leatf_top
(
input wire 	sys_clk,



)










divider_2s divider_2s_inst
(
.	sys_clk	(),

.clk_1s		(),
.clk_1ms	(),
.clk_1us    ()
);















endmodule 